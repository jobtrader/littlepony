library verilog;
use verilog.vl_types.all;
entity counter_debounce_vlg_vec_tst is
end counter_debounce_vlg_vec_tst;
